magic
tech sky130l
timestamp 1671835323
<< ndiffusion >>
rect 8 22 13 23
rect 8 19 9 22
rect 12 19 13 22
rect 8 13 13 19
rect 15 13 20 23
rect 22 17 27 23
rect 22 14 23 17
rect 26 14 27 17
rect 22 13 27 14
rect 33 17 38 23
rect 33 14 34 17
rect 37 14 38 17
rect 33 13 38 14
rect 40 17 45 23
rect 51 22 56 23
rect 51 19 52 22
rect 55 19 56 22
rect 51 17 56 19
rect 58 22 65 23
rect 58 19 60 22
rect 63 19 65 22
rect 58 17 65 19
rect 40 14 41 17
rect 44 14 45 17
rect 40 13 45 14
rect 61 13 65 17
rect 67 17 72 23
rect 67 14 68 17
rect 71 14 72 17
rect 67 13 72 14
<< ndc >>
rect 9 19 12 22
rect 23 14 26 17
rect 34 14 37 17
rect 52 19 55 22
rect 60 19 63 22
rect 41 14 44 17
rect 68 14 71 17
<< ntransistor >>
rect 13 13 15 23
rect 20 13 22 23
rect 38 13 40 23
rect 56 17 58 23
rect 65 13 67 23
<< pdiffusion >>
rect 8 47 13 48
rect 8 44 9 47
rect 12 44 13 47
rect 8 41 13 44
rect 8 38 9 41
rect 12 38 13 41
rect 8 33 13 38
rect 15 41 19 48
rect 33 47 38 48
rect 33 44 34 47
rect 37 44 38 47
rect 33 41 38 44
rect 15 40 20 41
rect 15 37 16 40
rect 19 37 20 40
rect 15 33 20 37
rect 22 37 27 41
rect 22 34 23 37
rect 26 34 27 37
rect 22 33 27 34
rect 33 38 34 41
rect 37 38 38 41
rect 33 33 38 38
rect 40 47 45 48
rect 40 44 41 47
rect 44 44 45 47
rect 40 41 45 44
rect 40 38 41 41
rect 44 38 45 41
rect 40 33 45 38
rect 51 47 56 48
rect 51 44 52 47
rect 55 44 56 47
rect 51 41 56 44
rect 51 38 52 41
rect 55 38 56 41
rect 51 33 56 38
rect 58 33 65 48
rect 67 47 72 48
rect 67 44 68 47
rect 71 44 72 47
rect 67 41 72 44
rect 67 38 68 41
rect 71 38 72 41
rect 67 33 72 38
<< pdc >>
rect 9 44 12 47
rect 9 38 12 41
rect 34 44 37 47
rect 16 37 19 40
rect 23 34 26 37
rect 34 38 37 41
rect 41 44 44 47
rect 41 38 44 41
rect 52 44 55 47
rect 52 38 55 41
rect 68 44 71 47
rect 68 38 71 41
<< ptransistor >>
rect 13 33 15 48
rect 20 33 22 41
rect 38 33 40 48
rect 56 33 58 48
rect 65 33 67 48
<< polysilicon >>
rect 13 48 15 50
rect 38 48 40 50
rect 56 48 58 50
rect 65 48 67 50
rect 20 41 22 43
rect 13 30 15 33
rect 9 29 15 30
rect 9 26 10 29
rect 13 26 15 29
rect 9 25 15 26
rect 13 23 15 25
rect 20 30 22 33
rect 38 30 40 33
rect 56 30 58 33
rect 20 29 26 30
rect 20 26 22 29
rect 25 26 26 29
rect 20 25 26 26
rect 33 29 40 30
rect 33 26 34 29
rect 37 26 40 29
rect 33 25 40 26
rect 52 29 58 30
rect 52 26 53 29
rect 56 26 58 29
rect 52 25 58 26
rect 20 23 22 25
rect 38 23 40 25
rect 56 23 58 25
rect 65 23 67 33
rect 13 11 15 13
rect 20 10 22 13
rect 38 11 40 13
rect 56 10 58 17
rect 65 11 67 13
rect 20 9 25 10
rect 20 6 21 9
rect 24 6 25 9
rect 20 5 25 6
rect 53 9 58 10
rect 53 6 54 9
rect 57 6 58 9
rect 62 10 67 11
rect 62 7 63 10
rect 66 7 67 10
rect 62 6 67 7
rect 53 5 58 6
<< pc >>
rect 10 26 13 29
rect 22 26 25 29
rect 34 26 37 29
rect 53 26 56 29
rect 21 6 24 9
rect 54 6 57 9
rect 63 7 66 10
<< m1 >>
rect 42 51 45 57
rect 9 47 12 48
rect 9 41 12 44
rect 9 37 12 38
rect 16 40 19 49
rect 41 48 45 51
rect 34 47 37 48
rect 34 41 37 44
rect 34 37 37 38
rect 41 47 44 48
rect 41 41 44 44
rect 41 37 44 38
rect 52 47 55 48
rect 52 41 55 44
rect 52 37 55 38
rect 68 47 71 49
rect 68 41 71 44
rect 68 37 71 38
rect 16 36 19 37
rect 22 34 23 37
rect 26 34 31 37
rect 22 29 25 30
rect 9 26 10 29
rect 13 26 14 29
rect 28 29 31 34
rect 53 29 56 30
rect 28 26 34 29
rect 37 26 50 29
rect 22 25 25 26
rect 9 22 12 23
rect 47 22 50 26
rect 53 25 56 26
rect 60 22 63 23
rect 47 19 52 22
rect 55 19 56 22
rect 9 18 12 19
rect 60 18 63 19
rect 34 17 37 18
rect 22 14 23 17
rect 26 14 34 17
rect 34 13 37 14
rect 41 17 44 18
rect 41 13 44 14
rect 68 17 71 18
rect 68 13 71 14
rect 74 10 77 38
rect 21 9 24 10
rect 54 9 57 10
rect 24 6 54 7
rect 62 7 63 10
rect 66 7 67 10
rect 21 4 57 6
rect 21 2 24 4
rect 63 2 66 7
<< m2c >>
rect 16 49 19 52
rect 9 38 12 41
rect 68 49 71 52
rect 34 38 37 41
rect 41 38 44 41
rect 52 38 55 41
rect 74 38 77 41
rect 10 26 13 29
rect 22 26 25 29
rect 9 19 12 22
rect 53 26 56 29
rect 60 19 63 22
rect 41 14 44 17
rect 68 14 71 17
rect 34 10 37 13
rect 74 7 77 10
<< m2 >>
rect 15 52 20 53
rect 15 51 16 52
rect 4 49 16 51
rect 19 51 20 52
rect 67 52 72 53
rect 67 51 68 52
rect 19 49 68 51
rect 71 49 72 52
rect 15 48 20 49
rect 67 48 72 49
rect 8 41 13 42
rect 33 41 38 42
rect 8 38 9 41
rect 12 39 34 41
rect 12 38 13 39
rect 8 37 13 38
rect 33 38 34 39
rect 37 38 38 41
rect 33 37 38 38
rect 40 41 45 42
rect 40 38 41 41
rect 44 39 45 41
rect 51 41 56 42
rect 51 39 52 41
rect 44 38 52 39
rect 55 39 56 41
rect 73 41 78 42
rect 73 39 74 41
rect 55 38 74 39
rect 77 38 78 41
rect 40 37 78 38
rect 9 29 14 30
rect 4 27 10 29
rect 9 26 10 27
rect 13 26 14 29
rect 9 25 14 26
rect 21 29 26 30
rect 52 29 57 30
rect 21 26 22 29
rect 25 27 53 29
rect 25 26 26 27
rect 21 25 26 26
rect 52 26 53 27
rect 56 26 57 29
rect 52 25 57 26
rect 8 22 82 23
rect 8 19 9 22
rect 12 21 60 22
rect 12 19 13 21
rect 8 18 13 19
rect 59 19 60 21
rect 63 21 82 22
rect 63 19 64 21
rect 59 18 64 19
rect 40 17 45 18
rect 40 14 41 17
rect 44 15 45 17
rect 67 17 72 18
rect 67 15 68 17
rect 44 14 68 15
rect 71 14 72 17
rect 33 13 38 14
rect 40 13 72 14
rect 33 10 34 13
rect 37 11 38 13
rect 37 10 78 11
rect 33 9 74 10
rect 73 7 74 9
rect 77 7 78 10
rect 73 6 78 7
<< labels >>
rlabel space 0 -4 0 -4 3 WARNINGS
rlabel m2 16 53 16 53 5 EXTEND_Vdd_HERE
rlabel m2 72 39 72 39 1 Vdd
port 1 n
rlabel space 0 -8 0 -8 3 Router's_path_to_GND_is_blocked
rlabel m2 62 14 62 14 1 GND
port 2 n
rlabel m1 67 8 67 8 1 B
port 3 n
rlabel space 0 -12 0 -12 3 Router's_path_to_A_is_blocked
rlabel polysilicon 14 12 14 12 1 A
port 4 n
rlabel m2 57 11 57 11 1 S
port 5 n
rlabel m2 56 39 56 39 1 Y
port 6 n
rlabel m2 78 8 78 8 7 M2_ON_EDGE
rlabel m2c 75 8 75 8 1 M2_ON_EDGE
rlabel m2 74 7 74 7 1 M2_ON_EDGE
rlabel m2 74 8 74 8 1 M2_ON_EDGE
rlabel m2 38 11 38 11 1 M2_ON_EDGE
rlabel m2 38 12 38 12 1 M2_ON_EDGE
rlabel m2c 35 11 35 11 1 M2_ON_EDGE
rlabel m2 34 10 34 10 1 M2_ON_EDGE
rlabel m2 34 11 34 11 1 M2_ON_EDGE
rlabel m2 34 14 34 14 1 M2_ON_EDGE
<< end >>
